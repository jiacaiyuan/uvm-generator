`ifndef {{ module.upper() }}_ENV_PKG_SVH
`define {{ module.upper() }}_ENV_PKG_SVH

  `include "{{ module }}_env_config.sv"
  `include "{{ module }}_virtual_sequencer.sv"
  `include "{{ module }}_env_checker.sv"
  `include "{{ module }}_env.sv"

`endif