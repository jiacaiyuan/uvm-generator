`ifndef {{ module.upper() }}_COMMON_PKG_SVH
`define {{ module.upper() }}_COMMON_PKG_SVH

  `include "{{ module }}_type.sv"
  `include "{{ module }}_agent_config.sv"
  `include "{{ module }}_item.sv"

`endif